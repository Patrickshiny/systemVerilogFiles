package uvm_custom_pkg;
	import uvm_pkg::*;
	class uvm_custom_env extends uvm_env;
    endclass
endpackage
