module top_module(
    output logic zero
);
  assign zero = 0;
endmodule
